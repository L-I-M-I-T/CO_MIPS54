`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/07/14 23:46:11
// Design Name: 
// Module Name: MULT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MULT(
input [31:0] a,
input [31:0] b,
output [63:0] z
);

wire [63:0] a1;
wire [64:0] z1;

assign a1=(a[31]==0)?{32'b00000000000000000000000000000000,a}:{32'b11111111111111111111111111111111,a};
assign z1=((b[0]?a1:65'b0)+((b[1]==1)?(a1<<1):65'b0)+((b[2]==1)?(a1<<2):65'b0)+((b[3]==1)?(a1<<3):65'b0)+((b[4]==1)?(a1<<4):65'b0)+((b[5]==1)?(a1<<5):65'b0)+((b[6]==1)?(a1<<6):65'b0)+((b[7]==1)?(a1<<7):65'b0)+((b[8]==1)?(a1<<8):65'b0)+((b[9]==1)?(a1<<9):65'b0)+((b[10]==1)?(a1<<10):65'b0)+((b[11]==1)?(a1<<11):65'b0)+((b[12]==1)?(a1<<12):65'b0)+((b[13]==1)?(a1<<13):65'b0)+((b[14]==1)?(a1<<14):65'b0)+((b[15]==1)?(a1<<15):65'b0)+((b[16]==1)?(a1<<16):65'b0)+((b[17]==1)?(a1<<17):65'b0)+((b[18]==1)?(a1<<18):65'b0)+((b[19]==1)?(a1<<19):65'b0)+((b[20]==1)?(a1<<20):65'b0)+((b[21]==1)?(a1<<21):65'b0)+((b[22]==1)?(a1<<22):65'b0)+((b[23]==1)?(a1<<23):65'b0)+((b[24]==1)?(a1<<24):65'b0)+((b[25]==1)?(a1<<25):65'b0)+((b[26]==1)?(a1<<26):65'b0)+((b[27]==1)?(a1<<27):65'b0)+((b[28]==1)?(a1<<28):65'b0)+((b[29]==1)?(a1<<29):65'b0)+((b[30]==1)?(a1<<30):65'b0)-((b[31]==1)?a1<<31:65'b0));
assign z=z1[63:0];

endmodule
